`timescale 1ns / 1ps

/*

*/

module fig_08a_block_200(
	input all_bits_pending,
	input plot,
	input rpix,
	input ram_done,
	input pleq,
	input scr_md,
	
	output dump,
	output clrpnd,
	output ldpnd,
	output ldpix,
	output bpr );
	
	


endmodule
