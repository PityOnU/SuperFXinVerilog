`timescale 1ns / 1ps

/*


*/

module fig_04b_block_076_078(
	input clk,
	input enable,
	input data_in,
	input disable_l,
	input enable_h,
	input disable_h,
	input cchld,
	input pcen,
	input loopen,
	input reset,
	input rn15,
	output [15:0] x,
	output [15:0] y
    );


endmodule
